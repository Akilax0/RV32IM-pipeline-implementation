module alu_tb;


endmodule
