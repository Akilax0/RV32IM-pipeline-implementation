`include "./alu.v"
`include "./reg_file.v"

module cpu();
//================= STAGE 1 ==========================



//================= STAGE 2 ==========================
//================= STAGE 3 ==========================
//================= STAGE 4 ==========================
//================= STAGE 5 ==========================


endmodule
